

class test1 extends uvm_test;

endclass