
class driver1 extends uvm_driver;

endclass